package rob_pkg;

  `include "sys_defs.svh"
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "sequence_item.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "coverage.sv"
  `include "scoreboard.sv"
  `include "agent.sv"
  `include "env.sv"
  `include "base_seq.sv"
  `include "reset_seq.sv"
  `include "random_seq.sv"
  `include "test.sv"

endpackage : rob_pkg